module normalize_ff(
P,
P_normalized
);



endmodule
